/******************************filter module*************************************/
/*property:Interpolated FIR
/*fpass:40Hz
/*fstop:100Hz
/*FS:@7812.5Hz
/*Numerator:									binary:(*8192)					decimal:(*8192)
				0.056190570395043708					111001100							460
				0.057164981312558115					111010100							468
				0.058018058683830982					111011100							476
				0.058746166444177433					111100001							481
				0.059346193853615406					111100110							486
				0.059815572373094157					111101010							490
				0.060152289616208533					111101101							493
				0.060354900290602947					111101110							494
				0.060422534061737462					111110000							496
				0.060354900290602947					111101110							494
				0.060152289616208533					111101101							493
				0.059815572373094157					111101010							490
				0.059346193853615406					111100110							486
				0.058746166444177433					111100001							481
				0.058018058683830982					111011100							476
				0.057164981312558115					111010100							468
				0.056190570395043708					111001100							460
/***********************************end******************************************/
module adc_fir (fir_clk,rst,adc_indata,adc_outdata);

input wire fir_clk,rst;
input wire [15:0] adc_indata;
output wire [15:0] adc_outdata;

reg [15:0] r0,r1,r2,r3,r4,r5,r6,r7,r8,r9,r10,r11,r12,r13,r14,r15,r16;
always @ (posedge fir_clk,negedge rst)
	begin
		if (!rst)
			begin
				r0<=16'd0;r1<=16'd0;r2<=16'd0;r3<=16'd0;r4<=16'd0;r5<=16'd0;r6<=16'd0;r7<=16'd0;r8<=16'd0;r9<=16'd0;r10<=16'd0;r11<=16'd0;r12<=16'd0;r13<=16'd0;r14<=16'd0;r15<=16'd0;r16<=16'd0;
			end 
		else 
			begin
				r0<=adc_indata;
				r1<=r0;
				r2<=r1;
				r3<=r2;
				r4<=r3;
				r5<=r4;
				r6<=r5;
				r7<=r6;
				r8<=r7;
				r9<=r8;
				r10<=r9;
				r11<=r10;
				r12<=r11;
				r13<=r12;
				r14<=r13;
				r15<=r14;
//				r16<=r15;
			end  
	end
//wire [27:0] c0,c1,c2,c3,c4,c5,c6,c7,c8,c9,c10,c11,c12,c13,c14,c15,c16;
//assign c0={{r0,2'd0}+{r0,3'd0}+{r0,6'd0}+{r0,7'd0}+{r0,8'd0}};
//assign c1={{r1,2'd0}+{r1,4'd0}+{r1,6'd0}+{r1,7'd0}+{r1,8'd0}};
//assign c2={{r2,2'd0}+{r2,3'd0}+{r2,4'd0}+{r2,6'd0}+{r2,7'd0}+{r2,8'd0}};
//assign c3={r3+{r3,5'd0}+{r3,6'd0}+{r3,7'd0}+{r3,8'd0}};
//assign c4={{r4,1'd0}+{r4,2'd0}+{r4,5'd0}+{r4,6'd0}+{r4,7'd0}+{r4,8'd0}};
//assign c5={{r5,1'd0}+{r5,3'd0}+{r5,5'd0}+{r5,6'd0}+{r5,7'd0}+{r5,8'd0}};
//assign c6={r6+{r6,2'd0}+{r6,3'd0}+{r6,5'd0}+{r6,6'd0}+{r6,7'd0}+{r6,8'd0}};
//assign c7={{r7,1'd0}+{r7,2'd0}+{r7,3'd0}+{r7,5'd0}+{r7,6'd0}+{r7,7'd0}+{r7,8'd0}};
//assign c8={{r8,4'd0}+{r8,5'd0}+{r8,6'd0}+{r8,7'd0}+{r8,8'd0}};
//assign c9={{r9,1'd0}+{r9,2'd0}+{r9,3'd0}+{r9,5'd0}+{r9,6'd0}+{r9,7'd0}+{r9,8'd0}};
//assign c10={r10+{r10,2'd0}+{r10,3'd0}+{r10,5'd0}+{r10,6'd0}+{r10,7'd0}+{r10,8'd0}};
//assign c11={{r11,1'd0}+{r11,3'd0}+{r11,5'd0}+{r11,6'd0}+{r11,7'd0}+{r11,8'd0}};
//assign c12={{r12,1'd0}+{r12,2'd0}+{r12,5'd0}+{r12,6'd0}+{r12,7'd0}+{r12,8'd0}};
//assign c13={r13+{r13,5'd0}+{r13,6'd0}+{r13,7'd0}+{r13,8'd0}};
//assign c14={{r14,2'd0}+{r14,3'd0}+{r14,4'd0}+{r14,6'd0}+{r14,7'd0}+{r14,8'd0}};
//assign c15={{r15,2'd0}+{r15,4'd0}+{r15,6'd0}+{r15,7'd0}+{r15,8'd0}};
//assign c16={{r16,2'd0}+{r16,3'd0}+{r16,6'd0}+{r16,7'd0}+{r16,8'd0}};

//assign c0=r0*9'd460;
//assign c1=r1*9'd468;
//assign c2=r2*9'd476;
//assign c3=r3*9'd481;
//assign c4=r4*9'd486;
//assign c5=r5*9'd490;
//assign c6=r6*9'd493;
//assign c7=r7*9'd494;
//assign c8=r8*9'd496;
//assign c9=r9*9'd494;
//assign c10=r10*9'd493;
//assign c11=r11*9'd490;
//assign c12=r12*9'd486;
//assign c13=r13*9'd481;
//assign c14=r14*9'd476;
//assign c15=r15*9'd468;
//assign c16=r16*9'd460;

//reg [28:0] sum;
//always @ (posedge fir_clk,negedge rst)
//	begin
//		if (!rst)
//			sum<=29'd0;
//		else
//			sum=c0+c1+c2+c3+c4+c5+c6+c7+c8+c9+c10+c11+c12+c13+c14+c15+c16;
//	end

wire [20:0] sum;
assign sum=r0+r1+r2+r3+r4+r5+r6+r7+r8+r9+r10+r11+r12+r13+r14+r15;

assign adc_outdata=sum[20:5];
	
endmodule  